
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:38:09 02/04/2012 
// Design Name: 
// Module Name:    ioTest 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: Testing IO board.
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ioTest (input  M_CLOCK,
					input  [3:0] btn,       // IO Board Pushbutton Switches 
					output reg [3:0] an, 	// IO Board Seven Segment Digits					
					output reg [7:0] seg,   // 7=dp, 6=g, 5=f,4=e, 3=d,2=c,1=b, 0=a
					output reg dp);         // Decimal point in the seven segment
					
					// active low
					
					
					IO_SSEG = 4'b1110;
					
					case



endmodule
	